library verilog;
use verilog.vl_types.all;
entity calc_if is
    port(
        clk             : in     vl_logic
    );
end calc_if;
