`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x0+qddVU5c2vjHYytU2y85FwN3W/fRKTvvtsQI/HbifJ/GfQIW0J8Vr3TgBp1ZXI
59gtgF5GrcVF4xr2iqiLV82GVznNjilhqRWPNcn4Uh9Ey1AtwaW1D4qEYUhO/Q/8
OMMYgZMDbE1aRC0EdW+7z5Dvm4qT1Yj9PfxY+rlN6HGv3cz/Igl/BvqW4fDGq1qo
OPduw2WcolGFnSdXtwK0pWwx/u1zGiv1EDNa0t0y5XKZ9PCgq7Ba6mbo+K10E2OB
G1qnoLoU4vQrmk6b/xVaz/idMMheJ6DU1W086pkZKzf+fe7py2P9MaDWSLX3LthM
nN5TZd+93gyM02tQhDjK92Id2MGnvHmAaCExMsgUcaDQgbgSiZP8qtFfJopwASTH
VgWj+SXbXtE9q3tK1hk3mcqgV5gei6BkDd0ONAtWgBCMEP6U0aZumzaRimHbD8wJ
kxC3B8doyZ7eOPhTGdGegN7FUNXChNEk7XV9XXhys7r1d96NJW+ucZJ02z56RVT5
/dcon7EnkAi/yDqxccaTZq7ngh3TninA6NDcnxarGmr02QCVL9QkkPMkjFOXhFL9
BHX2InF7lxF2sezkGYt5NOABA7jt+3++lLy6wDTMbUtsQpNitb+muB00N/LmrAFu
Fd6hnCc4i29VHsZSywJAM6xceMWpKygk3yAyLyJMnLcuuDYROXzTESW3wVfHTPde
j/B/VLSPRVLUtad9nFwL1i9X1x95bgzUMHEpLnk5fwsWe0u8JqUC6nKeEWyQhrqp
N/k3iUTZw4Wk7P51D/6syQuahj7y08XwbAfE4tKxshZq7mOgCMiQWU0fMhBXM4sz
jbMyiltNR8kS0H/yqazHqNxvdLBMqrKk8RXGzYUjjAkqd1IrQCs4ehUWmm9hnrQT
TC+Yrr/ecMTaBvAOkF2EZofdGz2zQkYrvbabdQD5w3eZb3tOerrQQyvsYh7D9GZt
kqkBvmuuIUltCY8gwxcGIRoebRdI8HJ7vVB4UybsXEERP6qE/H8RnpGcoHKjsHHV
cK5zsDeuisZQwYAn/NUKrxuDdpAD4mAvglgAJtQgJbe69xngNXXF7TPe/NDdjkcC
qrXwyrxd1lpC4SM2UPYZE//e41ZaN+oSvSUk9vXPl9JlkRtF+gvuqbogU1TRZGDS
KS9+/3DwfHlaY3jarz9Wsnps0OQLbSb3EcAnT0D1dKojWqJHjHwqAhIL8kmSFNZK
Pax7XdRd5Du16+V2Yzovw7ZpPNPotMwJr14rDCIQpaDv5cx7ggtclXoJpXyWz7Lv
Le+vueIVmrRTQi4tCyA9iwUoLySgv0t8/gvkJ5eAiN/IujaDEypXcsY4aknTxn05
wZ62DK2oicDYNsaF/ixxll813QyaO6AW6BgiDZag2uERpQe8w8EhqgV3mkZjri6l
0DiqvVq4Vt1dw+48B67lQ1nTN5j5hOv8ozcJr8zmZQjTMvuYi0w1Dhw95YlnpXvm
lhrrKnx9SnDFHzlMc4KMdjAM0psKWzQoB3jA89wB8+IdN2a94pRz/T4lixphJ83N
KYtK1RXiys6hoLzWj/0kAmSp2S4QF82olzknkaemT1i0++AbCNurS40dbmRR7w7/
+jVGGrBjphCei9WzmupTu24hrHZJ0s/7dNk+tfgiui1y0bfI7J6FTW9vjWEcQvFq
81yf+NQmEkZVIS9T+MLJYa9O72VxEZDrR5oUK7nIItF4FtnWSF9lM2IKQvW939eR
I0pY3Oj58gSypYgrMma1HstbwJPXdo6ObPntZ1qmXcPiyqqi57Zlfw8akeFJvPzv
4ZJx77Vmskn79VaHYHKP1Mx91dovudSzd6ERwNM8rDthLYPN0zFFPrmd8F91hi4y
Uxm9HnwPX2Xz8t+iAblyjLSRunZZdcpQ5sHEHz56XJAeuZUiXQ7oa5EY/7pHlMlp
5D1HYgvKHW7tyx3MQrQ4bK1+34eMFyJe4BgwCpuQp6O0OsOM74CR5bAjG9M3CLL7
tC+HKe4mkgSHfX0DY4DnXGSnE/SezmibrkLe1qnnZMCv9sxC1yfej97rveePueII
fGIAsCsprOJXXKxgvSHEYKtf2/whsJTTmHzljEKNXB4QIHBaIzjIOyYVcAfow4FY
KPcNlYOdUeeWxgdkvyA4tvTmjlBHPHNY7xwGE4CMaObTeBZgxeFpGLkYO+7rJQKJ
710pqzFVBRzEzkRPQP3Vk2R3FIGzBIWrFdmd/LSGdGVgJDMz4aF+Q75ZNnluVJXM
gF/uhbY6e/K+z4sxQ/1ViD/4Ge18vVPYMOT4gs0YidAYw+9VA5mcQxsF/CoNm+4I
PPLKsUGM+uf8kpuH74CUW3PqxsbfXomOWVUEwJ7JWNNfEZvHWJWsenfPRLzvRoI/
iki1mzydPZTTvzzERbZEt0Al3161kqrZPY+Ovwdo6NnJAlGtps472l0ouPe83J7R
HfSB4IhqPS3q+mvjHiYPniLD8jJw8vh7XHvLySLu52JhfRE4f+7DRV0K3AlZMKBb
N6CJSY00Pvp4SxpJLxqlogsNwjPe0Oj8WUGjvFq8rHMm9fY9PqM1NEIQdStYEo7W
beH2jCMk4cf733p0asHrT1Kpsl5Gis1Q11sNH0usbvmEi5b1QOZNPlmoXnTamICC
R4c1YnlAKPfpqpXEjNJS9saCk9TFprtrMRZ1OmLi8x1nRM1deoEb9a2UgQVYzUCq
ZdPZMhIjFnGzYrR27m2AIoCK2RxbYtdOX8/ROdBgeZXLBTtQUy1ImUDOJOsn6/Er
SIE4fGVaOeqfmkM6Zv94Qt392TH14UEcJ06s36ZyvcPy6MH4TpXXt6EQ/tl49ugw
p7u44xyZzJsgqNOD/5jvrpydlTtiiIorgiLbQ9N1G1wD/gxo4479Hb42cvRYF1U3
AjqSqVwIyZasaKLpPG8RbGaBLRinZpl57t0rsPuryE3R8yzO8AlJbfAYmhARuGPN
+oc4poBqG4QUL/TyPiLobzMl0ZkdQA9E/ualP1QOvb3/4/LEfjnX2N+t0oe/Rls4
uGKQS26R7PdJ1PIKe87+Xb7SSahmxzyyYQPZ8NGbOVD3j0IE9YTOUJaEwpnMqhXh
FeYZcC7vGekXvB7i7zU1xQ==
`protect END_PROTECTED
