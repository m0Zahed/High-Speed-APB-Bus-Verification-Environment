library verilog;
use verilog.vl_types.all;
entity calc_if_sv_unit is
end calc_if_sv_unit;
