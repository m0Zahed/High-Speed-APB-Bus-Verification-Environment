`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2e0LKl2SBR1NkY47j92mRN11Qsk+CJHQZh2njQJsIjEdw9+mJ8nbl0GUxCa64623
uafkiyoCwTdfLJ6fpogNXIJboawgXfrm14/IzRJd3ACca8AEhbiQKuOmMk8M1yJ5
n/D8PsYjIXQ/s0uyeKBqE0HawmQgqw+mU67GJwtdjOlytJP0hHLxntfwtpQ2SnWn
Z+JEi3vURmFavlHvYTJGaArgISFFcXc00gPZLAbTnGw0i9Yj2gIezW3iXiHCZvuS
YlrHVIHgeLgUjbWrAF5r/jHxL3/lNpC2fehDiNjpkiFKHXtjnbFbVmZbC7aBOFNg
qK+uh6TcmOrZVHE+obzqTqVqMGHXmKc/Xxv1CmMkKAGWg9fcPLAARW56aHA19aPj
JAGQVG2C3AVOlboBeHy5qdGYK8Uab/SZew0hSmZ7ZvOibG961PlQb0tN/OEVRko3
2S7BbninwbMPYjFTYemYONWNKZ2ACV5LFn6yIQuX6dXbxzzxT0tATG1JbGU1XAlv
`protect END_PROTECTED
