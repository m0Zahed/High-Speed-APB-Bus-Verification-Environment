`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hfNOXd8YJHccJkyrf+5P+wdaHAIJbxJt4cD9jDFMD7bmQ/WBHUiMdTEOdDRnCC1y
DHaovAuOwdQhhBR/C9UMsGII06mlatmtwTbXYKrVKDLsP87JSHUTtQq6BNhrg82P
hTmt8hZITVyJ/Kf8z0sc7G9Wlu5Yd9/ZXLP7LVSxmTQadUjUO52XJOzN95XL3CaN
3TsReshTBZhDrAWNGBynHx+Z8Rkk9UomMPlhMrB1fNsSCBCOGKwu9Q+2kY44cSDY
SSnU5cMhUGRM4e8L2tsLMMGguFJgvZvT0raujOTwqx9Sg1gc5M0qRzGyw08oLzfi
okHu48Uka13IelH21kCG1zrv9DElOcwOTjh7DmBpG0kzenjygexj/LgkKD2CJ0SC
vgTFRDxpGbi0pJdGa6FUaqlnCVAU+lamfaDTDG6Ec4WPrOZPWr4ZS8GRynb8BWlF
vhc/7DykoGUU7owUEdhIRgUhP1fQmP59H6lF9oJ5aBdEC98kkyl3ZRaMP8/1r+Cf
ZZbS/ySY6GwYQe1XC6be6wwOYpoVO2CzndLX1cMvj2EECcld1PtXCmdn4RMeqd9k
fgOLoIRC/+6imsMsV0+gRZuEdp7luzbYgLI0f0GcB9vjnPbWcJNBLfbQpkETqkmv
`protect END_PROTECTED
