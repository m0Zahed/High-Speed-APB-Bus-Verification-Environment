`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8nSpMTT/EVjbG5QLHpmYkfEGAfqWQDvU6FmeNbnoCnYIdZKPwsU2iVMJyehlIesg
4Q+ScgKpAuOyRaHuIuiWuy8/U11DGnrLPXcPp9whNA1GmKpQ1Hg7NLtacIo4uztF
4RMhX+FNGBIMH6Z/Tua7Mg2zjQv3GH3ZzefrjZeAet26FQfvx8SLLyPBbVKv8kU6
I024wvUqKRkcN8odG3hlyYscP/WtzdPhMerQzNEhjwJ9p9fbOPHUhcuuDc7cGSPM
A/sYc2cro5Mhd7+Y+ZTdJvZ0FLZAjsXdGwsbhL4GJpxpU2kyEoRCyVAZS7LMQEo5
GkUBFFm0C6jtXxPHbcqS8COr5nnxYah4/LJYlsqFrsW7oK9AOzULG4hLZcrXaxZD
Ck7TDImgQv6Iwwz0jTo8Zekev+fdpXEd9JZFoukL8GxKajHJ+si0dD7zYPWC6UjM
8okM28L7GVIlM+G0q5WWKJsgUcveB8Jq3+z7SkyVzEn+tvMud7xgsykCUSDpumUT
KDHwiNFSM3UPuR1HnzAd4QDhsny3KEPw49EdEX9wJp11K206Ws8fg/9PolaKPJ+5
jj6WRjywx4pKidMVx5pIQHifwG5N0CfcaUL5pX2cnSPfRhlBwCyOTA3x/snQVUvu
Ulj2J+qsSH8I9tNNzP582yPg6q/ySXxl7bwRWoDZpNIfLFxjyg5cIfhaZTB2elsd
RBA/EAlKnQgQsKG9b1fzexXxiCFsqpyE4zxckczxjsLud9EHEPdNKltEtO+IzYkJ
c4RW1jSz1luw23dZ7AKH/akpbRdRkynLggGS02jWbYl1qydNjXRzLnIED932g16n
5GO9zaLnBMP9oLXBmKHum1XNtB+JL7DvkbphZRSyOeg=
`protect END_PROTECTED
