`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NaRqYuW8nu9Ym0mgKDN/G+x/BbzzWxkg913KEVMEaiODvZtr6/gWbdFod4EXtSAp
72aaoAI/0VvUnptIa4WStL3mQfT+W0dN5QOKA9+BkxNKQOBnjkTS2RQSVDcrJ3GA
BPmzKixTCXFFVU6eF7mbcGq2YrZdRp0+WtQvz6+jz/yBghCJZFuaUV9PNNT/c7iR
Ohr/qOvv3OGoQJ7ZU3p4f1oQqVr7OfPWq5//axmw5MrB3Xf87+7DdChQJ7x9CxYG
rlMFId4WNdUSmh0vbpjQT0rk99K4LoqD2DGkBdMAY+/67+DWUC5EaKoVxgw0aHWj
2FvAOsdRAKqQNQfXL0NgGfldm4LfLf6nhDO6Ub1hj0NPwzDgqXpfEsvUOlNNSMA2
gy6/pSRxikJuz3ZgjvxOF5VuxxUMqIEILfaFhKjLGUZ1p3v13UFifwU3xxUOj8wl
mDusIZ8ZnA3p3jictol0DYJQEnq1AUxN7E5g2GAgVUmDZ4pqe2baqGkqvltAtdKr
U/XNUtidolyPylA8i3wOf5svptkzj3IuWU8ihzyBcHWV/Hdt1JhZp+nAnKi2MBvw
UQRgZ+sOHUie+kuSvIZUeWfnLBgk9eHAnWiTWXbMbfyjf6Z24kwcpOai7blD5MuC
/fL7hQXpIO2VRQosE3ms05Yms9eXRfW8+FLvj3QFIanFd/GqZvBr1sfU+w6w3eOv
AbSQjQkvnwlMFzMuQ0oC18DPNraXp5w3Uc1gP1Fm5KGkqcBSzl9at9xQj+p7mbJp
vHyUJCTqSKkVgU6kc2K98027x+N5hsmiD8vc8UqVvRfdOPp2IWRa4hkhnZ8C1Y9j
64JbF23dy5Mqtk8CbPJy4SSKFRMgmD+2irRp0RblXveYW9RGaG+Vlmsvk3hrn3pY
8EnUfFS3yg9MzELOoXYaYJWlT+/zhLWBIjVshwNQCQLFvHslsH33qh4HwuYkFiIO
XUl7bBxwbCCBVdqYtLoG9T3Hpb44Yn1tVa5AN2sTTyh3AolAA1yniCfM7NoO/WNs
FMfuL6dVKOa7SrBjmA05TY/LgvkZnuggoGJ7VexiVfTz0BGT+5AnjPWSZaxSaWwY
fSm4oCQQec7IbrBZpu/jFqpBbQhCrUU1gplCJ/+bpN3lqHJV1EJVFtFEWMyE4QQ8
eP2YFl4d1IbNrv/+aWhIkVae1H9wJGYkaI7sjXtpxH4isTQgic52ojD0wTH8mXvS
HHzd51W8i17C7+5T3LQoEMy8CWB2qSU4k/PJP9w5QBKJ43rFmoAzgFIGlyQJA6NW
6l8o9k9EJGLJ+PVeN4qCxnGvoTmPvRmwJyRQOjIqkc/KPgirgAn5wKabj+qefDBr
GF3rfOYv19sWtSYw4mgyMMZeZ0yk4reKrlfN2jrGPDkjH3E7r0FvS02OG8mOXPet
QESsUB7SFZ6nNuKpzjN/fhuPVaBBlvNRtxRvNQDJT4+HsbKJ6HP8pPgB6b5gFppH
i0cCkG+XZAyxBoRVnG0nGhK/mRHKOBVN7C5mEykE41jw1Q5sxY1MIRaUTtD6AM3W
MLHwry27FXpw+UcloegY3Ng1X1rTnUO9iL1SaIob72mRnhMSrO5pfjP9JoAEHTYP
OcnwSRoGFXipfJ1dlAQsGOry9hNpwFUZAPn8Lv2F7Kpow7s/mpSBBT8/ZzL+IeLi
R7ICdrGCFUwM1o3di/jKvlyLM4ChSq4SWUYhk1DgVRW3XPNkKN/TMgAwIdjruJDN
`protect END_PROTECTED
