`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
e3vY2qNKd3tmYU/vf8OGc95lINGxOuzbCgCPyIUpxdEA1ytMvoS9htUCY04yROg9
yxm7yKZ1Za9iJdw553Udc3z8CgssXicGpzJ0+oKAJ+P4SNGJ+zgaRePntSGrDXlV
P2aQYbS24Bk3/omeZeygFBlSd/42UG3N8fjiT91ck3qtHYiJPdTNAXSzkw8ayDLE
RUI+jYyfy7ZTW3uT04rgaWqW+gP9T6nUEUgQ0EOtEuToIfFwmRg1LQBo+aABY3wk
H/rcaC2baO/UdNpgzJoXDgF7G0futOzbLyEbNZKvCAv879ZsdE5PA2LtnC3tLTLp
y3RXcYeMOZwnpjbez7Iu2n5YW9ex7ha0Te2bdP3ZuaHNqeE3BZ/WSTHu2X8ucVK+
0m0d2zKC/maOPbZYT4f7nMCmqNkGoJQbUTN0+4jwIXPwFJrdPFAYQurtQUvNKFZX
mO3gvVzkbbnZ0/Yn0LW8EqOlwIAM0oqNOHXqRvwAzUjl99dfVAcDe+ekCltZNJG8
UNI/LROpvCWEqYDKtiliUg/5qFGdjvjhwNfWqrppM/n3EJzygzMIHwyunTCCmhz1
wVteyrbE0g4MCqZrb4WaaRIxIhR67g49NjIDlZDtIrF6UKODo8DIsKOOoFd7F7w7
RYZtjJZ8pXUZUl3Hs0gBnkhiN08nReAdFNJhwAbfhA+m2tA1+TDvCdKZNPcxp6gz
4U9UtH/RLix1awYk2zQFA9LMuiyL+nrM2kS3hT1v9UWY39INmrAuxJh8ZHBhYnr4
ON2YAENrgCRIVGvrdl5CIqKmbKzYEzL2LMVuDv6izWtc45VP2r63a+S7ff5mSN5T
BaYvIsGZACMOTBz0ZJwKOdp6H2GfJnbhmcEdh3Q1fy/PCHAxZgVY4UtoH3WQFV1D
JTYNoNQfeevroOh4mLY3ZWwHz5xse1Dz1VSaGGOgGEKFnFNdK6KqD+RT7gs7PBYk
2YFOmMZjHvBsziLL/574gQbJGRPEINiFUhXfQCWrAuEEt3bV899y1EZ1rnSLgw4T
VrxBx8T4Nf53xR6VC6QUU5y3UqilgsInH9K6gi8VW1F2cAtKnf+n5XEShEaYNxrH
1Z13vQQPZ7IyEiWMXoAzr/roZRkSfsB5EVLVIEwbpKNVIzlndRxzMiflqIpDl3jf
5vnZAkjzeneOibX/eMEGnoUyQBO4/mLTe5hQyKoohxY+LOq6uaeejgrGZAmg8kcb
YlTFACbOzD7IhUM8+UC9VjJFe84SM/bwQATUnVca4MgQ397jL/Br0Bmgdk3PM7mh
f+XZ0TLAyjpGRhtF1Idf3W3jDE2iWUkwAYmdWUqhKwU=
`protect END_PROTECTED
