`ifndef __INFO__
`define __INFO__
class info;
    virtual function void display() 
      $display("Implement display function!"); 
    endfunction: display 
endclass : info
`endif
