`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NgI+xbm7K72lDkMXa6nCSntS45aDQZmXlkpbJMJh2xsYF2u4lC56BamdTK4SWyC1
FbyCkOPT5tcq1zwxsyKllyh5z45N9LuwOyAePiU8/73G0skguWtZx1CN9u2JPfCq
YL4mgeYtyXvuCfNPrxdvSdMRCNpswVxACb7Kbfk56cOzZ/PbxiTPr7s3lek71isD
M/j4NPhpu2Hj4hpr+zAonDqdQtb3T5q7Ama+cnx4wDRPc/UJNuTimVNaHTs0A796
MeunIN65M7hOexKbA5xJ7fP8cTiZEAegMKl5inlNSmuFCcjUfZRjc8ieuZEXFDFt
k2fED2vZcx2nlEhxvAfoiDJnZllxGlSiIN2S3j2ROm3C+cybJWKtyov1tFQZvnxM
68Y5dJ3QTAe1/a1ipgvMFQBw10xhGFUkiFX1cGbXAxydKTwPpk73eYlxyin7cF36
Db4Mx84Uh4Kq5dGfuV6XOzcwQZ8L4nMrxtPPmDPY6Xq8cE6kWrZYKDc0iHigUHoE
VjVKQVRGDc1yc/3iZTpNznCqeLJeeknrNWzbJshr3n0Xvw170IplDUc/Q9EjdnGI
E5dUPFUm0aIr9BAZwL6rlNPfOvNHVAZ10Dn8JuZumWagVO2YO5NSPnvlgCQ3omrF
v7kBfURtGXtJtvigVQw/g+GYi0Bv+UNTid+ACIFrQaRq7GcFzlrAaTRwJ1gGbSMs
fkWAJAkaMPRo9Z3W7Y1oN3egLbXtyKIDOf76JVJ7kZHQpet1T4K1pApZ70cBftfa
kj64d5G3bbJXnwqVb2ZI/MlidEKaTISAAmQZPWz1qLUM5MbQGie/yur3jB+/zt76
ZQy7XPMMgHsYhTTzd8mW7PDctG+wD8nlR2U365VFNRyRYDVOTQFaZ3aUyPiOwXRj
BzUAkPDkybZ5bLh9veBdvvi1K5WyCZ3v20KDblLK/YgJbFXdyFvqIVqZMiHs99qr
ZRBuyDVEuagg/QaU6GRfGbn3kydQcJTHFTqRqUWj19UdrHztkG4UMxrR4ZvX9JYN
0heUf/CqYqhuWBFDk89KTQ==
`protect END_PROTECTED
